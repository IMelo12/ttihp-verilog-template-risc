module tt_um_risc(
    input  wire [7:0] ui_in,    // Dedicated inputs
    output wire [7:0] uo_out,   // Kept as wire
    input  wire [7:0] uio_in,   // IOs: Input path
    output wire [7:0] uio_out,  // IOs: Output path
    output wire [7:0] uio_oe,   // IOs: Enable path (1=output)
    input  wire       ena,      // Enable signal
    input  wire       clk,      // Clock
    input  wire       rst_n     // Active-low reset
);

// Enable output on all uio pins
assign uio_oe = 8'hFF;

wire [7:0] risc_output;
wire input_we = ui_in[0];
wire [6:0] input_address = ui_in[7:1];
wire [7:0] input_data = uio_in;

(* dont_touch = "true" *) risc cpu(
    .clk(clk),
    .rst_n(rst_n),
    .inst_address(input_address),
    .inst_data(input_data),
    .inst_we(input_we),
    .memory_out(risc_output)
);

// Drive risc output to uio and uo
assign uio_out = risc_output;

// Example control: override output if ui_in == 8'b00000001 and ena is high
assign uo_out = (!rst_n)            ? 8'b0 :
                (ena && ui_in == 8'b00000001) ? 8'b1 :
                risc_output;

endmodule
